`timescale 1ns / 1ps

module testbench;
  reg clk;
  reg rst;
  reg C1;
  wire clockout;
  main testbench(.clk(clk),.clockout(clockout),.rst(rst),.C1(C1));
  initial
   begin
     $dumpfile("testbench.vcd");
     $dumpvars(0,testbench);
     clk = 0;
     rst = 0;
     C1=1;
     #50
     rst = 1;
     #10
     rst = 0;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     rst = 1;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     rst=0;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     C1 = 0;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #10 clk = ~clk;
     #100
     $finish;
   end
      
endmodule
